/**
 * @Author: German Cano Quiveu <germancq>
 * @Date:   2019-03-01T15:43:26+01:00
 * @Email:  germancq@dte.us.es
 * @Filename: autotest_module.v
 * @Last modified by:   germancq
 * @Last modified time: 2019-03-01T15:48:59+01:00
 */
module autotest_module(

  );

  fsm_autotest fsm_isnt(

  );


  sdspihost sdspi_inst(

  );

endmodule
