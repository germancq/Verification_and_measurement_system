/**
 * @ Author: German Cano Quiveu, germancq
 * @ Create Time: 2019-12-19 13:34:50
 * @ Modified by: Your name
 * @ Modified time: 2019-12-19 13:44:17
 * @ Description:
 */

package configuration;

    localparam N = 88;
    localparam DATA_WIDTH = 64;
    localparam c = 80;
    localparam r = 8;
    localparam R = 45;
    localparam lCounter_initial_state = 6'h05;
    localparam lCounter_feedback_coeff = 7'h61;

endpackage
