// Design: and gate
// Description: 
// Author: German Cano Quiveu <germancq@dte.us.es>
// Copyright Universidad de Sevilla, Spain
// Rev: 4, sep 2017

module and_gate(
	input a,
	input b,
	output c);

assign c = a & b;

endmodule
